`timescale 1ns / 1ps

module neural_network #(
    parameter INTEGER_BITS = 9,
    parameter FIXED_POINT_BITS = 4
)(
input        i_clk,
input i_reset,
input[INTEGER_BITS+FIXED_POINT_BITS-1:0] pool_output,
input pool_output_valid,
output reg[(INTEGER_BITS+FIXED_POINT_BITS)*2-1:0] neurons,
output reg output_valid
    );
    
    reg[INTEGER_BITS+FIXED_POINT_BITS-1:0] w1[5:0][5:0],w2[5:0][5:0], b1,b2, n1, n2;
    reg[3:0] row,col;
    reg[(INTEGER_BITS+FIXED_POINT_BITS)*2-1:0] temp1,temp2;
    
    initial begin
        w1[0][0] = 13'b0000000010000;
        w1[0][1] = 13'b0000000010000;
        w1[0][2] = 13'b0000000010000;
        w1[0][3] = 13'b0000000010000;
        w1[0][4] = 13'b0000000010000;
        w1[0][5] = 13'b0000000010000;
        w1[1][0] = 13'b0000000010000;
        w1[1][1] = 13'b0000000010000;
        w1[1][2] = 13'b0000000010000;
        w1[1][3] = 13'b0000000010000;
        w1[1][4] = 13'b0000000010000;
        w1[1][5] = 13'b0000000010000;
        w1[2][0] = 13'b0000000010000;
        w1[2][1] = 13'b0000000010000;
        w1[2][2] = 13'b0000000010000;
        w1[2][3] = 13'b0000000010000;
        w1[2][4] = 13'b0000000010000;
        w1[2][5] = 13'b0000000010000;
        w1[3][0] = 13'b0000000010000;
        w1[3][1] = 13'b0000000010000;
        w1[3][2] = 13'b0000000010000;
        w1[3][3] = 13'b0000000010000;
        w1[3][4] = 13'b0000000010000;
        w1[3][5] = 13'b0000000010000;
        w1[4][0] = 13'b0000000010000;
        w1[4][1] = 13'b0000000010000;
        w1[4][2] = 13'b0000000010000;
        w1[4][3] = 13'b0000000010000;
        w1[4][4] = 13'b0000000010000;
        w1[4][5] = 13'b0000000010000;
        w1[5][0] = 13'b0000000010000;
        w1[5][1] = 13'b0000000010000;
        w1[5][2] = 13'b0000000010000;
        w1[5][3] = 13'b0000000010000;
        w1[5][4] = 13'b0000000010000;
        w1[5][5] = 13'b0000000010000;
        
        w2[0][0] = 13'b0000000010000;
        w2[0][1] = 13'b0000000010000;
        w2[0][2] = 13'b0000000010000;
        w2[0][3] = 13'b0000000010000;
        w2[0][4] = 13'b0000000010000;
        w2[0][5] = 13'b0000000010000;
        w2[1][0] = 13'b0000000010000;
        w2[1][1] = 13'b0000000010000;
        w2[1][2] = 13'b0000000010000;
        w2[1][3] = 13'b0000000010000;
        w2[1][4] = 13'b0000000010000;
        w2[1][5] = 13'b0000000010000;
        w2[2][0] = 13'b0000000010000;
        w2[2][1] = 13'b0000000010000;
        w2[2][2] = 13'b0000000010000;
        w2[2][3] = 13'b0000000010000;
        w2[2][4] = 13'b0000000010000;
        w2[2][5] = 13'b0000000010000;
        w2[3][0] = 13'b0000000010000;
        w2[3][1] = 13'b0000000010000;
        w2[3][2] = 13'b0000000010000;
        w2[3][3] = 13'b0000000010000;
        w2[3][4] = 13'b0000000010000;
        w2[3][5] = 13'b0000000010000;
        w2[4][0] = 13'b0000000010000;
        w2[4][1] = 13'b0000000010000;
        w2[4][2] = 13'b0000000010000;
        w2[4][3] = 13'b0000000010000;
        w2[4][4] = 13'b0000000010000;
        w2[4][5] = 13'b0000000010000;
        w2[5][0] = 13'b0000000010000;
        w2[5][1] = 13'b0000000010000;
        w2[5][2] = 13'b0000000010000;
        w2[5][3] = 13'b0000000010000;
        w2[5][4] = 13'b0000000010000;
        w2[5][5] = 13'b0000000010000;
         
        b1 = 13'b0000000010000;
        b2 = 13'b0000000010000;
    end
    
    always @(posedge i_reset) begin
        row = 0;
        col=0;
        n1 = b1;
        n2 = b2;
        output_valid = 0; 
        neurons=0;
     end
     
     always @(posedge i_clk) begin
        if(pool_output_valid) begin
            if (!(row==6 && col==6)) begin
            temp1 = n1 + w1[row][col]*pool_output;
            n1 = temp1[INTEGER_BITS+2*FIXED_POINT_BITS-1:FIXED_POINT_BITS-1];
            temp2 = n2 + w2[row][col]*pool_output;
            n2 = temp2[INTEGER_BITS+2*FIXED_POINT_BITS-1:FIXED_POINT_BITS-1];
            end
            
            if (row<6) row = row+1;
            
            else if(col<6) begin
                row=0;
                col = col+1;                
            end
            
            else begin
                output_valid = 1;
                neurons = {n1,n2};
            end
        end
     end
    
    
endmodule
